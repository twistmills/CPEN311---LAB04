module decode(
	input clk,

	
);



endmodule